`ifndef DEFINES_HEADER_SVH
`define DEFINES_HEADER_SVH

`define EXCEPTION_WIDTH   4
`define ALU_CONTROL_WIDTH 7
`define XLEN              32

localparam logic [6:0]
    OPCODE_RESET    = 7'b000_0000,
    OPCODE_LOAD     = 7'b000_0011,
    OPCODE_FENCE    = 7'b000_1111,
    OPCODE_I_TYPE   = 7'b001_0011,
    OPCODE_AUIPC    = 7'b001_0111,
    OPCODE_S_TYPE   = 7'b010_0011,
    OPCODE_R_TYPE   = 7'b011_0011,
    OPCODE_LUI      = 7'b011_0111,
    OPCODE_B_TYPE   = 7'b110_0011,
    OPCODE_JALR     = 7'b110_0111,
    OPCODE_J_TYPE   = 7'b110_1111,
    OPCODE_SYSTEM   = 7'b111_0011,
    OPCODE_LOAD_FP  = 7'b000_0111,
    OPCODE_STORE_FP = 7'b010_0111,
    OPCODE_MADD     = 7'b100_0011,
    OPCODE_MSUB     = 7'b100_0111,
    OPCODE_NMSUB    = 7'b100_1011,
    OPCODE_NMADD    = 7'b100_1111,
    OPCODE_FP       = 7'b101_0011;

localparam logic [`ALU_CONTROL_WIDTH-1:0] 
    ALU_ADD       = 'b0000000,
    ALU_SUB       = 'b0000001,
    ALU_AND       = 'b0000010,
    ALU_OR        = 'b0000011,
    ALU_XOR       = 'b0000100,
    ALU_SLT       = 'b0000101,
    ALU_SLTU      = 'b0000110,
    ALU_SLL       = 'b0000111,
    ALU_SRL       = 'b0001000,
    ALU_SRA       = 'b0001001,
    ALU_PASS      = 'b0001010,
    
    ALU_MUL       = 'b0001011,
    ALU_MULH      = 'b0001100, 
    ALU_MULHSU    = 'b0001101, 
    ALU_MULHU     = 'b0001110, 
    ALU_DIV       = 'b0001111, 
    ALU_DIVU      = 'b0010000, 
    ALU_REM       = 'b0010001, 
    ALU_REMU      = 'b0010010, 
    
    ALU_ANDN      = 'b0010011, 
    ALU_ORN       = 'b0010100, 
    ALU_XNOR      = 'b0010101, 
    ALU_BCLR      = 'b0010110, 
    ALU_BEXT      = 'b0010111, 
    ALU_BINV      = 'b0011000, 
    ALU_BSET      = 'b0011001, 
    ALU_CLMUL     = 'b0011010, 
    ALU_CLMULH    = 'b0011011, 
    ALU_CLMULR    = 'b0011100, 
    ALU_MAX       = 'b0011101, 
    ALU_MAXU      = 'b0011110, 
    ALU_MIN       = 'b0011111, 
    ALU_MINU      = 'b0100000, 
    ALU_ROL       = 'b0100001, 
    ALU_ROR       = 'b0100010, 
    ALU_SH1ADD    = 'b0100011, 
    ALU_SH2ADD    = 'b0100100, 
    ALU_SH3ADD    = 'b0100101, 
    ALU_ZEXT_H    = 'b0100110, 
    ALU_CLZ       = 'b0101100, 
    ALU_CPOP      = 'b0101101, 
    ALU_CTZ       = 'b0101110, 
    ALU_ORC_B     = 'b0101111, 
    ALU_REV8      = 'b0110000, 
    ALU_SEXT_B    = 'b0110001, 
    ALU_SEXT_H    = 'b0110010,
    
    ALU_FLW       = 'b0110011,
    ALU_FSW       = 'b0110100,
    ALU_FMADD     = 'b0110101,
    ALU_FMSUB     = 'b0110110,
    ALU_FNMSUB    = 'b0110111,
    ALU_FNMADD    = 'b0111000,
    ALU_FADD      = 'b0111001,
    ALU_FSUB      = 'b0111010,
    ALU_FMUL      = 'b0111011,
    ALU_FDIV      = 'b0111100,
    ALU_FSQRT     = 'b0111101,
    ALU_FSGNJ     = 'b0111110,
    ALU_FSGNJN    = 'b0111111,
    ALU_FSGNJX    = 'b1000000,
    ALU_FMIN      = 'b1000001,
    ALU_FMAX      = 'b1000010,
    ALU_FCVTWS    = 'b1000011,
    ALU_FCVTWUS   = 'b1000100,
    ALU_FMVXW     = 'b1000101,
    ALU_FEQ       = 'b1000110,
    ALU_FLT       = 'b1000111,
    ALU_FLE       = 'b1001000,
    ALU_FCLASS    = 'b1001001,
    ALU_FCVTSW    = 'b1001010,
    ALU_FCVTSWU   = 'b1001011,
    ALU_FMVWX     = 'b1001100;

`endif // DEFINES_HEADER_SVH